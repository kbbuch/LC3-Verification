`ifndef PROTECT_PARAM
`define PROTECT_PARAM

parameter ADDX = 4'b0001;
parameter ANDX = 4'b0101;
parameter NOTX = 4'b1001;
parameter LDX =  4'b0010;
parameter LDRX = 4'b0110;
parameter LDIX = 4'b1010;
parameter LEAX = 4'b1110;
parameter STX =  4'b0011;
parameter STRX = 4'b0111;
parameter STIX = 4'b1011;
parameter BRX =  4'b0000;
parameter JMPX = 4'b1100;


`endif
